class {name} extends uvm_sequence_item;
    `uvm_object_utils({name})
    
    
  
    function new(string name = "{name}");
        super.new(name);
    endfunction
 
endclass : {name}